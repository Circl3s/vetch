module main

import getters as get

fn main() {
	print(get.user())
	print(get.host())
	print(get.uptime())
	print(get.os())
	print(get.version())
	print(get.term())
	print(get.shell())
	print(get.divider())
	print(get.cpu())
	print(get.gpu())
	print(get.memory())
	print(get.divider())
	print(get.colors())
}
